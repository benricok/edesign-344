* TIP41C NPN ho�drywingtransistor (TO220-pakkie)
.model TIP41C NPN(Is=457.5f Xti=3 Eg=1.11 Vaf=50 Bf=65 Ise=1.346p Ne=1.34
+          Ikf=3.296 Nc=.5961 Xtb=2.2 Br=7.639 Isc=604.1f Nc=2.168
+          Ikr=8.131m Rc=91.29m Cjc=278.7p Mjc=.385 Vjc=.75 Fc=.5 Cje=433p
+          Mje=.5 Vje=.75 Tr=1.412u Tf=37.34n Itf=35.68 Xtf=1.163 Vtf=10 Rb=.1)